// ------------------------------------------------------------------------------
//  POM employs sigma coordinates, which are bottom-following coordinates that map the vertical coordinate from
//  the vertical coordinate from -H < z < eta onto -1 < sigma_POM < 0, where z is -depth below ref level (not sea surface)
//  H > 0 is the static variable h(x,y) (in grid file) loaded into wdepth0
//  eta is dynamic variable elb(x,y) (in physics file) )
//  nz is number of faces vertically so that the number of wet cells is nz-1 vertically. 
//  Cell-centered arrays like t (temperature) are padded with an arbitrary value in last 
//  element iz=35 (surface cell at iz=1)
//  netCDF variable w(x,y,z) refers to vertical faces (not cell centers), so w(x,y,1) ~ 0 at sea surface and w(x,y,nz=35) = 0 at the sea bed.
//  Currently load these fields (in native units/conventions, c-declaration index order):
//     float elb(y, x)    = "surface elevation in external mode at -dt"  units = "metre" ;     staggering  = (east_e, north_e)
//     float u(z, y, x)   = "x-velocity"                                 units = "metre/sec" ; staggering  = (east_u, north_u, zz) 
//     float v(z, y, x)   = "y-velocity"                                 units = "metre/sec" ; staggering  = (east_v, north_v, zz) 
//     float w(z, y, x)   = "sigma-velocity"                             units = "metre/sec" ; staggering  = (east_e, north_e, z) 
//     float t(z, y, x)   = "potential temperature" ;                    units = "K" ;         staggering  = (east_e, north_e, zz) 
//     float s(z, y, x)   = "salinity x rho / rhoref" ;                  units = "PSS" ;       staggering  = (east_e, north_e, zz) 
//     float rho(z, y, x) = "(density-1000)/rhoref" ;                   units = "dimless"     staggering  = (east_e, north_e, zz)
//     float kh(z, y, x)  = "vertical diffusivity" ;                     units = "m^2/sec";    staggering  = (east_e, north_e, zz) 
//     float aam(z, y, x) = "horizontal kinematic viscosity" ;           units = "metre^2/sec";staggering  = (east_e, north_e, zz) 
//  u(ix,iy,iz) in grid position (ix-0.5, iy    , iz)     (i.e. western  cell face)
//  v(ix,iy,iz) in grid position (ix    , iy-0.5, iz)     (i.e. southern cell face)
//  w(ix,iy,iz) in grid position (ix    , iy,     iz-0.5) (i.e. upper    cell face)
//  The boundary condition:  w( ix, iy, nz+0.5 ) = 0   is implicit 
// ------------------------------------------------------------------------------
netcdf hydrography_YYYY_MM_DD {
dimensions:
	z = 35 ;
	y = 125 ;
	x = 182 ;
variables:
	float elb(y, x) ;
		elb:long_name = "surface elevation in external mode at -dt" ;
		elb:units = "metre" ;
		elb:coordinates = "east_e north_e" ;
	float u(z, y, x) ;
		u:long_name = "x-velocity" ;
		u:units = "metre/sec" ;
		u:coordinates = "east_u north_u zz" ;
	float v(z, y, x) ;
		v:long_name = "y-velocity" ;
		v:units = "metre/sec" ;
		v:coordinates = "east_v north_v zz" ;
	float w(z, y, x) ;
		w:long_name = "sigma-velocity" ;
		w:units = "metre/sec" ;
		w:coordinates = "east_e north_e zz" ;
	float t(z, y, x) ;
		t:long_name = "potential temperature" ;
		t:units = "K" ;
		t:coordinates = "east_e north_e zz" ;
	float s(z, y, x) ;
		s:long_name = "salinity x rho / rhoref" ;
		s:units = "PSS" ;
		s:coordinates = "east_e north_e zz" ;
	float rho(z, y, x) ;
		rho:long_name = "(density-1000)/rhoref" ;
		rho:units = "dimensionless" ;
		rho:coordinates = "east_e north_e zz" ;
	float kh(z, y, x) ;
		kh:long_name = "vertical diffusivity" ;
		kh:units = "metre^2/sec" ;
		kh:coordinates = "east_e north_e zz" ;
	float aam(z, y, x) ;
		aam:long_name = "horizontal kinematic viscosity" ;
		aam:units = "metre^2/sec" ;
		aam:coordinates = "east_e north_e zz" ;

// global attributes:
		:title = "black_sea" ;
		:description = "restart file" ;
}
